class i_sequencer extends uvm_sequencer #(seq_item );

    `uvm_component_utils(i_sequencer)

    function new(string name ,uvm_component parent);
        super.new(name,parent);
    endfunction 
    
endclass 